module dknf(
    input x1, x2, x3,
    output f4
);
    assign f4 = ~x1;  // ???????????? ??????? f4 = ~x1
endmodule
