library verilog;
use verilog.vl_types.all;
entity ddnf is
    port(
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        f4              : out    vl_logic
    );
end ddnf;
